    Library ieee;
    USE ieee.std_logic_vector.all;
    
    ENTITY MyEntity is
        port(
            clk : in std_logic;
            rst : in std_logic
        );
    end MyEntity;
